library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity resid_tb is
end entity;

architecture test of resid_tb is

component resid is
	generic (WIDTH_IN : integer := 128
	);
	port(	
	    hxRES	:	in  std_logic_vector(2*WIDTH_IN-1 downto 0);
		xMAC	:	in  std_logic_vector(3*WIDTH_IN-1 downto 0);
		EK	    :	in  std_logic_vector(4*WIDTH_IN-1 downto 0);
		res_id	:	out std_logic_vector(2*WIDTH_IN-1 downto 0);
		clk	    :	in  std_logic;
		reset	:	in  std_logic		
	);
end component;

CONSTANT WIDTH_IN : integer := 128;

CONSTANT clk_period : time := 1 ns;

Signal xEK :  std_logic_vector(4*WIDTH_IN-1 downto 0) := (4*WIDTH_IN-1 downto 0 => '0');
Signal xxMAC :  std_logic_vector(3*WIDTH_IN-1 downto 0) := (3*WIDTH_IN-1 downto 0 => '0');
Signal xhxRES :  std_logic_vector(2*WIDTH_IN-1 downto 0) := (2*WIDTH_IN-1 downto 0 => '0');
Signal res_id :  std_logic_vector(2*WIDTH_IN-1 downto 0) := (2*WIDTH_IN-1 downto 0 => '0');


Signal clk : std_logic := '0';
Signal reset_t : std_logic := '0';

Begin
	Aresid: resid 
		generic map(WIDTH_IN => WIDTH_IN)
		port map(	hxRES		=>	xhxRES,
				xMAC		=>	xxMAC,
				EK		=>	xEK,
				res_id		=>	res_id,
				clk		=>	clk,
				reset		=>	reset_t
		);
-- process for clock
clk_process : Process
Begin
	clk <= '0';
	wait for clk_period/2;
	clk <= '1';
	wait for clk_period/2;
end process;

stim_process: process
Begin

	reset_t <= '1';
	wait for 1 * clk_period;
	reset_t <= '0';
	wait for 1 * clk_period;
	
	xhxRES <= "0001110010111111111101111101001000110010101111001111001100001111110100010100000011100100110101010110110111010100011101101111101110010001001111100111010110111111011011101011000001001110100111000001011000101001001101001110000010010010001010111001110011110101";
	xxMAC <= "001011011001110111100001001001100001111010100101100101001110001001111110111110111110100101000011101011111011001101110011000101010000000000000011001011100011000100101001011111011100010000000101011010001110001110001110101110001000101000000110000000101100100101010001110000000110010111010110010100111100101110001110110001111001101110110111011110111110001011010001001000110111100000010100";
	xEK <= "01111100101100011010101000001101100010101110100100101010111000010001011011001110101001101101010010100001001110011000101010010011000111110000011001001100111101100000110101011011001110101000110101000011010010101101100101010010011010011101011011110000011101110101001010010011000011110011110001101100110010010010100000000000111100001011100100111101011111111010011111110000011100101010010000000101000111011001011111011111001111100111011001111000000110001101010000000111010101111000001001000110010100001111011000000101";
	
	wait for 100 * clk_period;

	wait;

end process;

end;

